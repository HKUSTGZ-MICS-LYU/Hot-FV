//Following code is from line 1
module b14(datao, wr, reset, clock, rd, addr, datai);

    input                clock;
    input                reset;
    input         [30:0] datai;
    output        [19:0] addr;
    output        [30:0] datao;
    output               rd;
    output               wr;
    reg  B = 1'b0;
    reg  [30:0] IR = 31'b0;
    reg  [19:0] addr = 20'b0;
    wire   cf;
    wire   clock;
    reg  [1:0]  d = 2'b0;
    wire  [30:0] datai;
    reg  [30:0] datao = 31'b0;
    wire  [2:0] df;
    wire  [3:0] ff;
    reg  [30:0] m = 31'b0;
    wire  [1:0] mf;
    reg  rd = 1'b0;
    reg  [30:0] reg0 = 31'b0;
    reg  [30:0] reg1 = 31'b0;
    reg  [30:0] reg2 = 31'b0;
    reg  [30:0] reg3 = 31'b0;
    wire   reset;
    reg  [30:0] rx = 31'b0;
    wire  [1:0] s;
    reg  state = 1'b0;
    reg  [30:0] t = 31'b0;
    wire  [19:0] tail;
    reg  wr = 1'b0;
    reg [999:0] coverage0 = 1000'b0;

    assign mf = IR[28:27];
  //assertion( mf = Extract(28, 27, IR)) 0
    assign df = IR[26:24];
  //assertion( df = Extract(26, 24, IR)) 1
    assign ff = IR[22:19];
  //assertion( ff = Extract(22, 19, IR)) 2
    assign cf = IR[23];
  //assertion( cf = Extract(23, 23, IR)) 3
    assign tail = IR[19:0];
  //assertion( tail = Extract(19, 0, IR)) 4
    assign s = IR[30:29];
  //assertion( s = Extract(30, 29, IR)) 5
    //Following code is from line 44
        always @(posedge clock) begin
            if ((reset == 1'b1))
                begin
                    coverage0[6] = 1;  //assertion( 1 == reset = True) 6
                    IR <= 31'h00000000;  //assertion( IR = 0) 8
                    d <= 2'h0;  //assertion( d = 0) 9
                    rx <= 31'h00000000;  //assertion( rx = 0) 10
                    m <= 31'h00000000;  //assertion( m = 0) 11
                    B <= 1'b0;  //assertion( B = 0) 12
                    reg0 <= 31'h00000000;  //assertion( reg0 = 0) 13
                    reg1 <= 31'h00000000;  //assertion( reg1 = 0) 14
                    reg2 <= 31'h00000000;  //assertion( reg2 = 0) 15
                    reg3 <= 31'h00000000;  //assertion( reg3 = 0) 16
                    addr <= 20'h00000;  //assertion( addr = 0) 17
                    rd <= 1'b0;  //assertion( rd = 0) 18
                    wr <= 1'b0;  //assertion( wr = 0) 19
                    datao <= 31'h00000000;  //assertion( datao = 0) 20
                    state <= 1'b0;  //assertion( state = 0) 21
                end
            else
                begin
                    coverage0[7] = 1;  //assertion( 1 == reset = False) 7
                    case (state)
                      1'b0:
                        begin
                            coverage0[22] = 1;  //assertion( 0 == state = True) 22
                            addr <= reg3[19:0];  //assertion( addr = Extract(19, 0, reg3)) 23
                            rd <= 1'b1;  //assertion( rd = 1) 24
                            IR <= datai;  //assertion( IR = datai) 25
                            state <= 1'b1;  //assertion( state = 1) 26
                            case (datai[30:29])
                              2'h0:
                                begin
                                    coverage0[27] = 1;  //assertion( 0 == Extract(30, 29, datai) = True) 27
                                    rx <= reg0;  //assertion( rx = reg0) 28
                                end
                              2'h1:
                                begin
                                    coverage0[29] = 1;  //assertion( 1 == Extract(30, 29, datai) = True) 29
                                    rx <= reg1;  //assertion( rx = reg1) 30
                                end
                              2'h2:
                                begin
                                    coverage0[31] = 1;  //assertion( 2 == Extract(30, 29, datai) = True) 31
                                    rx <= reg2;  //assertion( rx = reg2) 32
                                end
                              2'h3:
                                begin
                                    coverage0[33] = 1;  //assertion( 3 == Extract(30, 29, datai) = True) 33
                                    rx <= reg3;  //assertion( rx = reg3) 34
                                end
                            endcase
                        end
                      1'b1:
                        begin
                            coverage0[35] = 1;  //assertion( 1 == state = True) 35
                            case (cf)
                              1'b1:
                                begin
                                    coverage0[36] = 1;  //assertion( 1 == cf = True) 36
                                    case (mf)
                                      2'h0:
                                        begin
                                            coverage0[37] = 1;  //assertion( 0 == mf = True) 37
                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 38
                                        end
                                      2'h1:
                                        begin
                                            coverage0[39] = 1;  //assertion( 1 == mf = True) 39
                                            m = datai;  //assertion( m = datai) 40
                                            addr <= tail;  //assertion( addr = tail) 41
                                            rd <= 1'b1;  //assertion( rd = 1) 42
                                        end
                                      2'h2:
                                        begin
                                            coverage0[43] = 1;  //assertion( 2 == mf = True) 43
                                            addr <= (tail + reg1[19:0]);  //assertion( addr = tail + Extract(19, 0, reg1)) 44
                                            rd <= 1'b1;  //assertion( rd = 1) 45
                                            m = datai;  //assertion( m = datai) 46
                                        end
                                      2'h3:
                                        begin
                                            coverage0[47] = 1;  //assertion( 3 == mf = True) 47
                                            addr <= (tail + reg2[19:0]);  //assertion( addr = tail + Extract(19, 0, reg2)) 48
                                            rd <= 1'b1;  //assertion( rd = 1) 49
                                            m = datai;  //assertion( m = datai) 50
                                        end
                                    endcase
                                    case (ff)
                                      4'h0:
                                        begin
                                            coverage0[51] = 1;  //assertion( 0 == ff = True) 51
                                            if ((rx < m))
                                                begin
                                                    coverage0[52] = 1;  //assertion( ULT(rx, m) = True) 52
                                                    B <= 1'b1;  //assertion( B = 1) 54
                                                end
                                            else
                                                begin
                                                    coverage0[53] = 1;  //assertion( ULT(rx, m) = False) 53
                                                    B <= 1'b0;  //assertion( B = 0) 55
                                                end
                                        end
                                      4'h1:
                                        begin
                                            coverage0[56] = 1;  //assertion( 1 == ff = True) 56
                                            if ((rx >= m))
                                                begin
                                                    coverage0[57] = 1;  //assertion( UGE(rx, m) = True) 57
                                                    B <= 1'b1;  //assertion( B = 1) 59
                                                end
                                            else
                                                begin
                                                    coverage0[58] = 1;  //assertion( UGE(rx, m) = False) 58
                                                    B <= 1'b0;  //assertion( B = 0) 60
                                                end
                                        end
                                      4'h2:
                                        begin
                                            coverage0[61] = 1;  //assertion( 2 == ff = True) 61
                                            if ((rx == m))
                                                begin
                                                    coverage0[62] = 1;  //assertion( rx == m = True) 62
                                                    B <= 1'b1;  //assertion( B = 1) 64
                                                end
                                            else
                                                begin
                                                    coverage0[63] = 1;  //assertion( rx == m = False) 63
                                                    B <= 1'b0;  //assertion( B = 0) 65
                                                end
                                        end
                                      4'h3:
                                        begin
                                            coverage0[66] = 1;  //assertion( 3 == ff = True) 66
                                            if ((rx != m))
                                                begin
                                                    coverage0[67] = 1;  //assertion( rx != m = True) 67
                                                    B <= 1'b1;  //assertion( B = 1) 69
                                                end
                                            else
                                                begin
                                                    coverage0[68] = 1;  //assertion( rx != m = False) 68
                                                    B <= 1'b0;  //assertion( B = 0) 70
                                                end
                                        end
                                      4'h4:
                                        begin
                                            coverage0[71] = 1;  //assertion( 4 == ff = True) 71
                                            if ((rx <= m))
                                                begin
                                                    coverage0[72] = 1;  //assertion( ULE(rx, m) = True) 72
                                                    B <= 1'b1;  //assertion( B = 1) 74
                                                end
                                            else
                                                begin
                                                    coverage0[73] = 1;  //assertion( ULE(rx, m) = False) 73
                                                    B <= 1'b0;  //assertion( B = 0) 75
                                                end
                                        end
                                      4'h5:
                                        begin
                                            coverage0[76] = 1;  //assertion( 5 == ff = True) 76
                                            if ((rx > m))
                                                begin
                                                    coverage0[77] = 1;  //assertion( UGT(rx, m) = True) 77
                                                    B <= 1'b1;  //assertion( B = 1) 79
                                                end
                                            else
                                                begin
                                                    coverage0[78] = 1;  //assertion( UGT(rx, m) = False) 78
                                                    B <= 1'b0;  //assertion( B = 0) 80
                                                end
                                        end
                                      4'h6:
                                        begin
                                            coverage0[81] = 1;  //assertion( 6 == ff = True) 81
                                            if ((rx > 31'h3fffffff))
                                                begin
                                                    coverage0[82] = 1;  //assertion( UGT(rx, 1073741823) = True) 82
                                                    rx = rx;  //assertion( rx = rx) 84
                                                end
                                            else
                                                    coverage0[83] = 1;  //assertion( UGT(rx, 1073741823) = False) 83
                                            if ((rx < m))
                                                begin
                                                    coverage0[85] = 1;  //assertion( ULT(rx, m) = True) 85
                                                    B <= 1'b1;  //assertion( B = 1) 87
                                                end
                                            else
                                                begin
                                                    coverage0[86] = 1;  //assertion( ULT(rx, m) = False) 86
                                                    B <= 1'b0;  //assertion( B = 0) 88
                                                end
                                        end
                                      4'h7:
                                        begin
                                            coverage0[89] = 1;  //assertion( 7 == ff = True) 89
                                            if ((rx > 31'h3fffffff))
                                                begin
                                                    coverage0[90] = 1;  //assertion( UGT(rx, 1073741823) = True) 90
                                                    rx = rx;  //assertion( rx = rx) 92
                                                end
                                            else
                                                    coverage0[91] = 1;  //assertion( UGT(rx, 1073741823) = False) 91
                                            if ((rx >= m))
                                                begin
                                                    coverage0[93] = 1;  //assertion( UGE(rx, m) = True) 93
                                                    B <= 1'b1;  //assertion( B = 1) 95
                                                end
                                            else
                                                begin
                                                    coverage0[94] = 1;  //assertion( UGE(rx, m) = False) 94
                                                    B <= 1'b0;  //assertion( B = 0) 96
                                                end
                                        end
                                      4'h8:
                                        begin
                                            coverage0[97] = 1;  //assertion( 8 == ff = True) 97
                                            if (((rx < m) || (B == 1'b1)))
                                                begin
                                                    coverage0[98] = 1;  //assertion( Or(If(ULT(rx, m) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = True) 98
                                                    B <= 1'b1;  //assertion( B = 1) 100
                                                end
                                            else
                                                begin
                                                    coverage0[99] = 1;  //assertion( Or(If(ULT(rx, m) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = False) 99
                                                    B <= 1'b0;  //assertion( B = 0) 101
                                                end
                                        end
                                      4'h9:
                                        begin
                                            coverage0[102] = 1;  //assertion( 9 == ff = True) 102
                                            if (((~(rx < m)) || (B == 1'b1)))
                                                begin
                                                    coverage0[103] = 1;  //assertion( Or(If(Not(ULT(rx, m) == True) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = True) 103
                                                    B <= 1'b1;  //assertion( B = 1) 105
                                                end
                                            else
                                                begin
                                                    coverage0[104] = 1;  //assertion( Or(If(Not(ULT(rx, m) == True) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = False) 104
                                                    B <= 1'b0;  //assertion( B = 0) 106
                                                end
                                        end
                                      4'ha:
                                        begin
                                            coverage0[107] = 1;  //assertion( 10 == ff = True) 107
                                            if (((rx == m) || (B == 1'b1)))
                                                begin
                                                    coverage0[108] = 1;  //assertion( Or(If((rx == m) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = True) 108
                                                    B <= 1'b1;  //assertion( B = 1) 110
                                                end
                                            else
                                                begin
                                                    coverage0[109] = 1;  //assertion( Or(If((rx == m) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = False) 109
                                                    B <= 1'b0;  //assertion( B = 0) 111
                                                end
                                        end
                                      4'hb:
                                        begin
                                            coverage0[112] = 1;  //assertion( 11 == ff = True) 112
                                            if (((~(rx == m)) || (B == 1'b1)))
                                                begin
                                                    coverage0[113] = 1;  //assertion( Or(If(Not((rx == m) == True) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = True) 113
                                                    B <= 1'b1;  //assertion( B = 1) 115
                                                end
                                            else
                                                begin
                                                    coverage0[114] = 1;  //assertion( Or(If(Not((rx == m) == True) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = False) 114
                                                    B <= 1'b0;  //assertion( B = 0) 116
                                                end
                                        end
                                      4'hc:
                                        begin
                                            coverage0[117] = 1;  //assertion( 12 == ff = True) 117
                                            if (((~(rx > m)) || (B == 1'b1)))
                                                begin
                                                    coverage0[118] = 1;  //assertion( Or(If(Not(UGT(rx, m) == True) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = True) 118
                                                    B <= 1'b1;  //assertion( B = 1) 120
                                                end
                                            else
                                                begin
                                                    coverage0[119] = 1;  //assertion( Or(If(Not(UGT(rx, m) == True) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = False) 119
                                                    B <= 1'b0;  //assertion( B = 0) 121
                                                end
                                        end
                                      4'hd:
                                        begin
                                            coverage0[122] = 1;  //assertion( 13 == ff = True) 122
                                            if (((rx > m) || (B == 1'b1)))
                                                begin
                                                    coverage0[123] = 1;  //assertion( Or(If(UGT(rx, m) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = True) 123
                                                    B <= 1'b1;  //assertion( B = 1) 125
                                                end
                                            else
                                                begin
                                                    coverage0[124] = 1;  //assertion( Or(If(UGT(rx, m) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = False) 124
                                                    B <= 1'b0;  //assertion( B = 0) 126
                                                end
                                        end
                                      4'he:
                                        begin
                                            coverage0[127] = 1;  //assertion( 14 == ff = True) 127
                                            if ((rx > 31'h3fffffff))
                                                begin
                                                    coverage0[128] = 1;  //assertion( UGT(rx, 1073741823) = True) 128
                                                    rx = rx;  //assertion( rx = rx) 130
                                                end
                                            else
                                                    coverage0[129] = 1;  //assertion( UGT(rx, 1073741823) = False) 129
                                            if (((rx < m) || (B == 1'b1)))
                                                begin
                                                    coverage0[131] = 1;  //assertion( Or(If(ULT(rx, m) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = True) 131
                                                    B <= 1'b1;  //assertion( B = 1) 133
                                                end
                                            else
                                                begin
                                                    coverage0[132] = 1;  //assertion( Or(If(ULT(rx, m) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = False) 132
                                                    B <= 1'b0;  //assertion( B = 0) 134
                                                end
                                        end
                                      4'hf:
                                        begin
                                            coverage0[135] = 1;  //assertion( 15 == ff = True) 135
                                            if ((rx > 31'h3fffffff))
                                                begin
                                                    coverage0[136] = 1;  //assertion( UGT(rx, 1073741823) = True) 136
                                                    rx = rx;  //assertion( rx = rx) 138
                                                end
                                            else
                                                    coverage0[137] = 1;  //assertion( UGT(rx, 1073741823) = False) 137
                                            if (((~(rx < m)) || (B == 1'b1)))
                                                begin
                                                    coverage0[139] = 1;  //assertion( Or(If(Not(ULT(rx, m) == True) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = True) 139
                                                    B <= 1'b1;  //assertion( B = 1) 141
                                                end
                                            else
                                                begin
                                                    coverage0[140] = 1;  //assertion( Or(If(Not(ULT(rx, m) == True) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) = False) 140
                                                    B <= 1'b0;  //assertion( B = 0) 142
                                                end
                                        end
                                    endcase
                                end
                              1'b0:
                                begin
                                    coverage0[143] = 1;  //assertion( 0 == cf = True) 143
                                    if ((df != 3'h7))
                                        begin
                                            coverage0[144] = 1;  //assertion( 7 != df = True) 144
                                            if ((((df == 3'h5) && (B == 1'b0)) || ((df == 3'h4) && (B == 1'b1))))
                                                begin
                                                    coverage0[146] = 1;  //assertion( Or(If(And(If((5 == df) == True, 1, 0) == 1, If((0 == B) == True, 1, 0) == 1) == True, 1, 0) == 1, If(And(If((4 == df) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) == True, 1, 0) == 1) = True) 146
                                                    d = 2'h3;  //assertion( d = 3) 148
                                                end
                                            else
                                                begin
                                                    coverage0[147] = 1;  //assertion( Or(If(And(If((5 == df) == True, 1, 0) == 1, If((0 == B) == True, 1, 0) == 1) == True, 1, 0) == 1, If(And(If((4 == df) == True, 1, 0) == 1, If((1 == B) == True, 1, 0) == 1) == True, 1, 0) == 1) = False) 147
                                                    d = df[1:0];  //assertion( d = Extract(1, 0, df)) 149
                                                end
                                            case (ff)
                                              4'h0:
                                                begin
                                                    coverage0[150] = 1;  //assertion( 0 == ff = True) 150
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[151] = 1;  //assertion( 0 == mf = True) 151
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 152
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[153] = 1;  //assertion( 1 == mf = True) 153
                                                            m = datai;  //assertion( m = datai) 154
                                                            addr <= tail;  //assertion( addr = tail) 155
                                                            rd <= 1'b1;  //assertion( rd = 1) 156
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[157] = 1;  //assertion( 2 == mf = True) 157
                                                            addr <= (tail + reg1[19:0]);  //assertion( addr = tail + Extract(19, 0, reg1)) 158
                                                            rd <= 1'b1;  //assertion( rd = 1) 159
                                                            m = datai;  //assertion( m = datai) 160
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[161] = 1;  //assertion( 3 == mf = True) 161
                                                            addr <= (tail + reg2[19:0]);  //assertion( addr = tail + Extract(19, 0, reg2)) 162
                                                            rd <= 1'b1;  //assertion( rd = 1) 163
                                                            m = datai;  //assertion( m = datai) 164
                                                        end
                                                    endcase
                                                    t = 31'h00000000;  //assertion( t = 0) 165
                                                    case (d)
                                                      2'h0:
                                                        begin
                                                            coverage0[166] = 1;  //assertion( 0 == d = True) 166
                                                            reg0 = (t - m);  //assertion( reg0 = t - m) 167
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[168] = 1;  //assertion( 1 == d = True) 168
                                                            reg1 = (t - m);  //assertion( reg1 = t - m) 169
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[170] = 1;  //assertion( 2 == d = True) 170
                                                            reg2 = (t - m);  //assertion( reg2 = t - m) 171
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[172] = 1;  //assertion( 3 == d = True) 172
                                                            reg3 = (t - m);  //assertion( reg3 = t - m) 173
                                                        end
                                                    endcase
                                                end
                                              4'h1:
                                                begin
                                                    coverage0[174] = 1;  //assertion( 1 == ff = True) 174
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[175] = 1;  //assertion( 0 == mf = True) 175
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 176
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[177] = 1;  //assertion( 1 == mf = True) 177
                                                            m = datai;  //assertion( m = datai) 178
                                                            addr <= tail;  //assertion( addr = tail) 179
                                                            rd <= 1'b1;  //assertion( rd = 1) 180
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[181] = 1;  //assertion( 2 == mf = True) 181
                                                            addr <= (tail + reg1[19:0]);  //assertion( addr = tail + Extract(19, 0, reg1)) 182
                                                            rd <= 1'b1;  //assertion( rd = 1) 183
                                                            m = datai;  //assertion( m = datai) 184
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[185] = 1;  //assertion( 3 == mf = True) 185
                                                            addr <= (tail + reg2[19:0]);  //assertion( addr = tail + Extract(19, 0, reg2)) 186
                                                            rd <= 1'b1;  //assertion( rd = 1) 187
                                                            m = datai;  //assertion( m = datai) 188
                                                        end
                                                    endcase
                                                    reg2 = reg3;  //assertion( reg2 = reg3) 189
                                                    reg3 = m;  //assertion( reg3 = m) 190
                                                end
                                              4'h2:
                                                begin
                                                    coverage0[191] = 1;  //assertion( 2 == ff = True) 191
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[192] = 1;  //assertion( 0 == mf = True) 192
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 193
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[194] = 1;  //assertion( 1 == mf = True) 194
                                                            m = datai;  //assertion( m = datai) 195
                                                            addr <= tail;  //assertion( addr = tail) 196
                                                            rd <= 1'b1;  //assertion( rd = 1) 197
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[198] = 1;  //assertion( 2 == mf = True) 198
                                                            addr <= (tail + reg1[19:0]);  //assertion( addr = tail + Extract(19, 0, reg1)) 199
                                                            rd <= 1'b1;  //assertion( rd = 1) 200
                                                            m = datai;  //assertion( m = datai) 201
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[202] = 1;  //assertion( 3 == mf = True) 202
                                                            addr <= (tail + reg2[19:0]);  //assertion( addr = tail + Extract(19, 0, reg2)) 203
                                                            rd <= 1'b1;  //assertion( rd = 1) 204
                                                            m = datai;  //assertion( m = datai) 205
                                                        end
                                                    endcase
                                                    case (d)
                                                      2'h0:
                                                        begin
                                                            coverage0[206] = 1;  //assertion( 0 == d = True) 206
                                                            reg0 = m;  //assertion( reg0 = m) 207
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[208] = 1;  //assertion( 1 == d = True) 208
                                                            reg1 = m;  //assertion( reg1 = m) 209
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[210] = 1;  //assertion( 2 == d = True) 210
                                                            reg2 = m;  //assertion( reg2 = m) 211
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[212] = 1;  //assertion( 3 == d = True) 212
                                                            reg3 = m;  //assertion( reg3 = m) 213
                                                        end
                                                    endcase
                                                end
                                              4'h3:
                                                begin
                                                    coverage0[214] = 1;  //assertion( 3 == ff = True) 214
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[215] = 1;  //assertion( 0 == mf = True) 215
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 216
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[217] = 1;  //assertion( 1 == mf = True) 217
                                                            m = datai;  //assertion( m = datai) 218
                                                            addr <= tail;  //assertion( addr = tail) 219
                                                            rd <= 1'b1;  //assertion( rd = 1) 220
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[221] = 1;  //assertion( 2 == mf = True) 221
                                                            addr <= (tail + reg1[19:0]);  //assertion( addr = tail + Extract(19, 0, reg1)) 222
                                                            rd <= 1'b1;  //assertion( rd = 1) 223
                                                            m = datai;  //assertion( m = datai) 224
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[225] = 1;  //assertion( 3 == mf = True) 225
                                                            addr <= (tail + reg2[19:0]);  //assertion( addr = tail + Extract(19, 0, reg2)) 226
                                                            rd <= 1'b1;  //assertion( rd = 1) 227
                                                            m = datai;  //assertion( m = datai) 228
                                                        end
                                                    endcase
                                                    case (d)
                                                      2'h0:
                                                        begin
                                                            coverage0[229] = 1;  //assertion( 0 == d = True) 229
                                                            reg0 = m;  //assertion( reg0 = m) 230
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[231] = 1;  //assertion( 1 == d = True) 231
                                                            reg1 = m;  //assertion( reg1 = m) 232
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[233] = 1;  //assertion( 2 == d = True) 233
                                                            reg2 = m;  //assertion( reg2 = m) 234
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[235] = 1;  //assertion( 3 == d = True) 235
                                                            reg3 = m;  //assertion( reg3 = m) 236
                                                        end
                                                    endcase
                                                end
                                              4'h4:
                                                begin
                                                    coverage0[237] = 1;  //assertion( 4 == ff = True) 237
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[238] = 1;  //assertion( 0 == mf = True) 238
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 239
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[240] = 1;  //assertion( 1 == mf = True) 240
                                                            m = datai;  //assertion( m = datai) 241
                                                            addr <= tail;  //assertion( addr = tail) 242
                                                            rd <= 1'b1;  //assertion( rd = 1) 243
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[244] = 1;  //assertion( 2 == mf = True) 244
                                                            addr <= (tail + reg1[19:0]);  //assertion( addr = tail + Extract(19, 0, reg1)) 245
                                                            rd <= 1'b1;  //assertion( rd = 1) 246
                                                            m = datai;  //assertion( m = datai) 247
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[248] = 1;  //assertion( 3 == mf = True) 248
                                                            addr <= (tail + reg2[19:0]);  //assertion( addr = tail + Extract(19, 0, reg2)) 249
                                                            rd <= 1'b1;  //assertion( rd = 1) 250
                                                            m = datai;  //assertion( m = datai) 251
                                                        end
                                                    endcase
                                                    case (d)
                                                      2'h0:
                                                        begin
                                                            coverage0[252] = 1;  //assertion( 0 == d = True) 252
                                                            reg0 = (rx + m);  //assertion( reg0 = rx + m) 253
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[254] = 1;  //assertion( 1 == d = True) 254
                                                            reg1 = (rx + m);  //assertion( reg1 = rx + m) 255
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[256] = 1;  //assertion( 2 == d = True) 256
                                                            reg2 = (rx + m);  //assertion( reg2 = rx + m) 257
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[258] = 1;  //assertion( 3 == d = True) 258
                                                            reg3 = (rx + m);  //assertion( reg3 = rx + m) 259
                                                        end
                                                    endcase
                                                end
                                              4'h5:
                                                begin
                                                    coverage0[260] = 1;  //assertion( 5 == ff = True) 260
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[261] = 1;  //assertion( 0 == mf = True) 261
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 262
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[263] = 1;  //assertion( 1 == mf = True) 263
                                                            m = datai;  //assertion( m = datai) 264
                                                            addr <= tail;  //assertion( addr = tail) 265
                                                            rd <= 1'b1;  //assertion( rd = 1) 266
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[267] = 1;  //assertion( 2 == mf = True) 267
                                                            addr <= (tail + reg1[19:0]);  //assertion( addr = tail + Extract(19, 0, reg1)) 268
                                                            rd <= 1'b1;  //assertion( rd = 1) 269
                                                            m = datai;  //assertion( m = datai) 270
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[271] = 1;  //assertion( 3 == mf = True) 271
                                                            addr <= (tail + reg2[19:0]);  //assertion( addr = tail + Extract(19, 0, reg2)) 272
                                                            rd <= 1'b1;  //assertion( rd = 1) 273
                                                            m = datai;  //assertion( m = datai) 274
                                                        end
                                                    endcase
                                                    case (d)
                                                      2'h0:
                                                        begin
                                                            coverage0[275] = 1;  //assertion( 0 == d = True) 275
                                                            reg0 = (rx + m);  //assertion( reg0 = rx + m) 276
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[277] = 1;  //assertion( 1 == d = True) 277
                                                            reg1 = (rx + m);  //assertion( reg1 = rx + m) 278
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[279] = 1;  //assertion( 2 == d = True) 279
                                                            reg2 = (rx + m);  //assertion( reg2 = rx + m) 280
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[281] = 1;  //assertion( 3 == d = True) 281
                                                            reg3 = (rx + m);  //assertion( reg3 = rx + m) 282
                                                        end
                                                    endcase
                                                end
                                              4'h6:
                                                begin
                                                    coverage0[283] = 1;  //assertion( 6 == ff = True) 283
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[284] = 1;  //assertion( 0 == mf = True) 284
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 285
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[286] = 1;  //assertion( 1 == mf = True) 286
                                                            m = datai;  //assertion( m = datai) 287
                                                            addr <= tail;  //assertion( addr = tail) 288
                                                            rd <= 1'b1;  //assertion( rd = 1) 289
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[290] = 1;  //assertion( 2 == mf = True) 290
                                                            addr <= (tail + reg1[19:0]);  //assertion( addr = tail + Extract(19, 0, reg1)) 291
                                                            rd <= 1'b1;  //assertion( rd = 1) 292
                                                            m = datai;  //assertion( m = datai) 293
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[294] = 1;  //assertion( 3 == mf = True) 294
                                                            addr <= (tail + reg2[19:0]);  //assertion( addr = tail + Extract(19, 0, reg2)) 295
                                                            rd <= 1'b1;  //assertion( rd = 1) 296
                                                            m = datai;  //assertion( m = datai) 297
                                                        end
                                                    endcase
                                                    case (d)
                                                      2'h0:
                                                        begin
                                                            coverage0[298] = 1;  //assertion( 0 == d = True) 298
                                                            reg0 = (rx - m);  //assertion( reg0 = rx - m) 299
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[300] = 1;  //assertion( 1 == d = True) 300
                                                            reg1 = (rx - m);  //assertion( reg1 = rx - m) 301
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[302] = 1;  //assertion( 2 == d = True) 302
                                                            reg2 = (rx - m);  //assertion( reg2 = rx - m) 303
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[304] = 1;  //assertion( 3 == d = True) 304
                                                            reg3 = (rx - m);  //assertion( reg3 = rx - m) 305
                                                        end
                                                    endcase
                                                end
                                              4'h7:
                                                begin
                                                    coverage0[306] = 1;  //assertion( 7 == ff = True) 306
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[307] = 1;  //assertion( 0 == mf = True) 307
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 308
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[309] = 1;  //assertion( 1 == mf = True) 309
                                                            m = datai;  //assertion( m = datai) 310
                                                            addr <= tail;  //assertion( addr = tail) 311
                                                            rd <= 1'b1;  //assertion( rd = 1) 312
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[313] = 1;  //assertion( 2 == mf = True) 313
                                                            addr <= (tail + reg1[19:0]);  //assertion( addr = tail + Extract(19, 0, reg1)) 314
                                                            rd <= 1'b1;  //assertion( rd = 1) 315
                                                            m = datai;  //assertion( m = datai) 316
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[317] = 1;  //assertion( 3 == mf = True) 317
                                                            addr <= (tail + reg2[19:0]);  //assertion( addr = tail + Extract(19, 0, reg2)) 318
                                                            rd <= 1'b1;  //assertion( rd = 1) 319
                                                            m = datai;  //assertion( m = datai) 320
                                                        end
                                                    endcase
                                                    case (d)
                                                      2'h0:
                                                        begin
                                                            coverage0[321] = 1;  //assertion( 0 == d = True) 321
                                                            reg0 = (rx - m);  //assertion( reg0 = rx - m) 322
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[323] = 1;  //assertion( 1 == d = True) 323
                                                            reg1 = (rx - m);  //assertion( reg1 = rx - m) 324
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[325] = 1;  //assertion( 2 == d = True) 325
                                                            reg2 = (rx - m);  //assertion( reg2 = rx - m) 326
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[327] = 1;  //assertion( 3 == d = True) 327
                                                            reg3 = (rx - m);  //assertion( reg3 = rx - m) 328
                                                        end
                                                    endcase
                                                end
                                              4'h8:
                                                begin
                                                    coverage0[329] = 1;  //assertion( 8 == ff = True) 329
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[330] = 1;  //assertion( 0 == mf = True) 330
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 331
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[332] = 1;  //assertion( 1 == mf = True) 332
                                                            m = datai;  //assertion( m = datai) 333
                                                            addr <= tail;  //assertion( addr = tail) 334
                                                            rd <= 1'b1;  //assertion( rd = 1) 335
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[336] = 1;  //assertion( 2 == mf = True) 336
                                                            addr <= (tail + reg1[19:0]);  //assertion( addr = tail + Extract(19, 0, reg1)) 337
                                                            rd <= 1'b1;  //assertion( rd = 1) 338
                                                            m = datai;  //assertion( m = datai) 339
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[340] = 1;  //assertion( 3 == mf = True) 340
                                                            addr <= (tail + reg2[19:0]);  //assertion( addr = tail + Extract(19, 0, reg2)) 341
                                                            rd <= 1'b1;  //assertion( rd = 1) 342
                                                            m = datai;  //assertion( m = datai) 343
                                                        end
                                                    endcase
                                                    case (d)
                                                      2'h0:
                                                        begin
                                                            coverage0[344] = 1;  //assertion( 0 == d = True) 344
                                                            reg0 = (rx + m);  //assertion( reg0 = rx + m) 345
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[346] = 1;  //assertion( 1 == d = True) 346
                                                            reg1 = (rx + m);  //assertion( reg1 = rx + m) 347
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[348] = 1;  //assertion( 2 == d = True) 348
                                                            reg2 = (rx + m);  //assertion( reg2 = rx + m) 349
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[350] = 1;  //assertion( 3 == d = True) 350
                                                            reg3 = (rx + m);  //assertion( reg3 = rx + m) 351
                                                        end
                                                    endcase
                                                end
                                              4'h9:
                                                begin
                                                    coverage0[352] = 1;  //assertion( 9 == ff = True) 352
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[353] = 1;  //assertion( 0 == mf = True) 353
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 354
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[355] = 1;  //assertion( 1 == mf = True) 355
                                                            m = datai;  //assertion( m = datai) 356
                                                            addr <= tail;  //assertion( addr = tail) 357
                                                            rd <= 1'b1;  //assertion( rd = 1) 358
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[359] = 1;  //assertion( 2 == mf = True) 359
                                                            addr <= (tail + reg1[19:0]);  //assertion( addr = tail + Extract(19, 0, reg1)) 360
                                                            rd <= 1'b1;  //assertion( rd = 1) 361
                                                            m = datai;  //assertion( m = datai) 362
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[363] = 1;  //assertion( 3 == mf = True) 363
                                                            addr <= (tail + reg2[19:0]);  //assertion( addr = tail + Extract(19, 0, reg2)) 364
                                                            rd <= 1'b1;  //assertion( rd = 1) 365
                                                            m = datai;  //assertion( m = datai) 366
                                                        end
                                                    endcase
                                                    case (d)
                                                      2'h0:
                                                        begin
                                                            coverage0[367] = 1;  //assertion( 0 == d = True) 367
                                                            reg0 = (rx - m);  //assertion( reg0 = rx - m) 368
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[369] = 1;  //assertion( 1 == d = True) 369
                                                            reg1 = (rx - m);  //assertion( reg1 = rx - m) 370
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[371] = 1;  //assertion( 2 == d = True) 371
                                                            reg2 = (rx - m);  //assertion( reg2 = rx - m) 372
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[373] = 1;  //assertion( 3 == d = True) 373
                                                            reg3 = (rx - m);  //assertion( reg3 = rx - m) 374
                                                        end
                                                    endcase
                                                end
                                              4'ha:
                                                begin
                                                    coverage0[375] = 1;  //assertion( 10 == ff = True) 375
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[376] = 1;  //assertion( 0 == mf = True) 376
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 377
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[378] = 1;  //assertion( 1 == mf = True) 378
                                                            m = datai;  //assertion( m = datai) 379
                                                            addr <= tail;  //assertion( addr = tail) 380
                                                            rd <= 1'b1;  //assertion( rd = 1) 381
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[382] = 1;  //assertion( 2 == mf = True) 382
                                                            addr <= (tail + reg1[19:0]);  //assertion( addr = tail + Extract(19, 0, reg1)) 383
                                                            rd <= 1'b1;  //assertion( rd = 1) 384
                                                            m = datai;  //assertion( m = datai) 385
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[386] = 1;  //assertion( 3 == mf = True) 386
                                                            addr <= (tail + reg2[19:0]);  //assertion( addr = tail + Extract(19, 0, reg2)) 387
                                                            rd <= 1'b1;  //assertion( rd = 1) 388
                                                            m = datai;  //assertion( m = datai) 389
                                                        end
                                                    endcase
                                                    case (d)
                                                      2'h0:
                                                        begin
                                                            coverage0[390] = 1;  //assertion( 0 == d = True) 390
                                                            reg0 = (rx + m);  //assertion( reg0 = rx + m) 391
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[392] = 1;  //assertion( 1 == d = True) 392
                                                            reg1 = (rx + m);  //assertion( reg1 = rx + m) 393
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[394] = 1;  //assertion( 2 == d = True) 394
                                                            reg2 = (rx + m);  //assertion( reg2 = rx + m) 395
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[396] = 1;  //assertion( 3 == d = True) 396
                                                            reg3 = (rx + m);  //assertion( reg3 = rx + m) 397
                                                        end
                                                    endcase
                                                end
                                              4'hb:
                                                begin
                                                    coverage0[398] = 1;  //assertion( 11 == ff = True) 398
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[399] = 1;  //assertion( 0 == mf = True) 399
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 400
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[401] = 1;  //assertion( 1 == mf = True) 401
                                                            m = datai;  //assertion( m = datai) 402
                                                            addr <= tail;  //assertion( addr = tail) 403
                                                            rd <= 1'b1;  //assertion( rd = 1) 404
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[405] = 1;  //assertion( 2 == mf = True) 405
                                                            addr <= (tail + reg1[19:0]);  //assertion( addr = tail + Extract(19, 0, reg1)) 406
                                                            rd <= 1'b1;  //assertion( rd = 1) 407
                                                            m = datai;  //assertion( m = datai) 408
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[409] = 1;  //assertion( 3 == mf = True) 409
                                                            addr <= (tail + reg2[19:0]);  //assertion( addr = tail + Extract(19, 0, reg2)) 410
                                                            rd <= 1'b1;  //assertion( rd = 1) 411
                                                            m = datai;  //assertion( m = datai) 412
                                                        end
                                                    endcase
                                                    case (d)
                                                      2'h0:
                                                        begin
                                                            coverage0[413] = 1;  //assertion( 0 == d = True) 413
                                                            reg0 = (rx - m);  //assertion( reg0 = rx - m) 414
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[415] = 1;  //assertion( 1 == d = True) 415
                                                            reg1 = (rx - m);  //assertion( reg1 = rx - m) 416
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[417] = 1;  //assertion( 2 == d = True) 417
                                                            reg2 = (rx - m);  //assertion( reg2 = rx - m) 418
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[419] = 1;  //assertion( 3 == d = True) 419
                                                            reg3 = (rx - m);  //assertion( reg3 = rx - m) 420
                                                        end
                                                    endcase
                                                end
                                              4'hc:
                                                begin
                                                    coverage0[421] = 1;  //assertion( 12 == ff = True) 421
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[422] = 1;  //assertion( 0 == mf = True) 422
                                                            t = {1'b0, rx[30:1]};  //assertion( t = Concat(0, Extract(30, 1, rx))) 423
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[424] = 1;  //assertion( 1 == mf = True) 424
                                                            t = {1'b0, ((B == 1'b1) ? 1'b0 : rx[30]), rx[29:1]};  //assertion( t = Concat(Concat(0, If((1 == B) == True, 0, Extract(30, 30, rx))), Extract(29, 1, rx))) 425
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[426] = 1;  //assertion( 2 == mf = True) 426
                                                            t = {rx[29:0], 1'b0};  //assertion( t = Concat(Extract(29, 0, rx), 0)) 427
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[428] = 1;  //assertion( 3 == mf = True) 428
                                                            t = {rx[29:0], 1'b0};  //assertion( t = Concat(Extract(29, 0, rx), 0)) 429
                                                            if ((t > 31'h3fffffff))
                                                                begin
                                                                    coverage0[430] = 1;  //assertion( UGT(t, 1073741823) = True) 430
                                                                    B <= 1'b1;  //assertion( B = 1) 432
                                                                end
                                                            else
                                                                begin
                                                                    coverage0[431] = 1;  //assertion( UGT(t, 1073741823) = False) 431
                                                                    B <= 1'b0;  //assertion( B = 0) 433
                                                                end
                                                        end
                                                    endcase
                                                    case (d)
                                                      2'h0:
                                                        begin
                                                            coverage0[434] = 1;  //assertion( 0 == d = True) 434
                                                            reg0 <= t;  //assertion( reg0 = t) 435
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[436] = 1;  //assertion( 1 == d = True) 436
                                                            reg1 <= t;  //assertion( reg1 = t) 437
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[438] = 1;  //assertion( 2 == d = True) 438
                                                            reg2 <= t;  //assertion( reg2 = t) 439
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[440] = 1;  //assertion( 3 == d = True) 440
                                                            reg3 <= t;  //assertion( reg3 = t) 441
                                                        end
                                                    endcase
                                                end
                                            endcase
                                        end
                                    else
                                        begin
                                            coverage0[145] = 1;  //assertion( 7 != df = False) 145
                                            if ((df == 3'h7))
                                                begin
                                                    coverage0[442] = 1;  //assertion( 7 == df = True) 442
                                                    case (mf)
                                                      2'h0:
                                                        begin
                                                            coverage0[444] = 1;  //assertion( 0 == mf = True) 444
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 445
                                                        end
                                                      2'h1:
                                                        begin
                                                            coverage0[446] = 1;  //assertion( 1 == mf = True) 446
                                                            m = {11'h000, tail};  //assertion( m = Concat(0, tail)) 447
                                                        end
                                                      2'h2:
                                                        begin
                                                            coverage0[448] = 1;  //assertion( 2 == mf = True) 448
                                                            m = (reg1 + {11'h000, tail});  //assertion( m = reg1 + Concat(0, tail)) 449
                                                        end
                                                      2'h3:
                                                        begin
                                                            coverage0[450] = 1;  //assertion( 3 == mf = True) 450
                                                            m = (reg2 + {11'h000, tail});  //assertion( m = reg2 + Concat(0, tail)) 451
                                                        end
                                                    endcase
                                                    addr <= m[19:0];  //assertion( addr = Extract(19, 0, m)) 452
                                                    wr <= 1'b1;  //assertion( wr = 1) 453
                                                    datao <= rx;  //assertion( datao = rx) 454
                                                end
                                            else
                                                    coverage0[443] = 1;  //assertion( 7 == df = False) 443
                                        end
                                end
                            endcase
                            state <= 1'b0;  //assertion( state = 0) 455
                        end
                    endcase
                end
        end
                            assert property (coverage0[6]==0);

                    assert property (coverage0[7]==0);

                            assert property (coverage0[22]==0);

                                    assert property (coverage0[27]==0);

                                    assert property (coverage0[29]==0);

                                    assert property (coverage0[31]==0);

                                    assert property (coverage0[33]==0);

                            assert property (coverage0[35]==0);

                                    assert property (coverage0[36]==0);

                                            assert property (coverage0[37]==0);

                                            assert property (coverage0[39]==0);

                                            assert property (coverage0[43]==0);

                                            assert property (coverage0[47]==0);

                                            assert property (coverage0[51]==0);

                                                    assert property (coverage0[52]==0);

                                                    assert property (coverage0[53]==0);

                                            assert property (coverage0[56]==0);

                                                    assert property (coverage0[57]==0);

                                                    assert property (coverage0[58]==0);

                                            assert property (coverage0[61]==0);

                                                    assert property (coverage0[62]==0);

                                                    assert property (coverage0[63]==0);

                                            assert property (coverage0[66]==0);

                                                    assert property (coverage0[67]==0);

                                                    assert property (coverage0[68]==0);

                                            assert property (coverage0[71]==0);

                                                    assert property (coverage0[72]==0);

                                                    assert property (coverage0[73]==0);

                                            assert property (coverage0[76]==0);

                                                    assert property (coverage0[77]==0);

                                                    assert property (coverage0[78]==0);

                                            assert property (coverage0[81]==0);

                                                    assert property (coverage0[82]==0);

                                                    assert property (coverage0[83]==0);

                                                    assert property (coverage0[85]==0);

                                                    assert property (coverage0[86]==0);

                                            assert property (coverage0[89]==0);

                                                    assert property (coverage0[90]==0);

                                                    assert property (coverage0[91]==0);

                                                    assert property (coverage0[93]==0);

                                                    assert property (coverage0[94]==0);

                                            assert property (coverage0[97]==0);

                                                    assert property (coverage0[98]==0);

                                                    assert property (coverage0[99]==0);

                                            assert property (coverage0[102]==0);

                                                    assert property (coverage0[103]==0);

                                                    assert property (coverage0[104]==0);

                                            assert property (coverage0[107]==0);

                                                    assert property (coverage0[108]==0);

                                                    assert property (coverage0[109]==0);

                                            assert property (coverage0[112]==0);

                                                    assert property (coverage0[113]==0);

                                                    assert property (coverage0[114]==0);

                                            assert property (coverage0[117]==0);

                                                    assert property (coverage0[118]==0);

                                                    assert property (coverage0[119]==0);

                                            assert property (coverage0[122]==0);

                                                    assert property (coverage0[123]==0);

                                                    assert property (coverage0[124]==0);

                                            assert property (coverage0[127]==0);

                                                    assert property (coverage0[128]==0);

                                                    assert property (coverage0[129]==0);

                                                    assert property (coverage0[131]==0);

                                                    assert property (coverage0[132]==0);

                                            assert property (coverage0[135]==0);

                                                    assert property (coverage0[136]==0);

                                                    assert property (coverage0[137]==0);

                                                    assert property (coverage0[139]==0);

                                                    assert property (coverage0[140]==0);

                                    assert property (coverage0[143]==0);

                                            assert property (coverage0[144]==0);

                                                    assert property (coverage0[146]==0);

                                                    assert property (coverage0[147]==0);

                                                    assert property (coverage0[150]==0);

                                                            assert property (coverage0[151]==0);

                                                            assert property (coverage0[153]==0);

                                                            assert property (coverage0[157]==0);

                                                            assert property (coverage0[161]==0);

                                                            assert property (coverage0[166]==0);

                                                            assert property (coverage0[168]==0);

                                                            assert property (coverage0[170]==0);

                                                            assert property (coverage0[172]==0);

                                                    assert property (coverage0[174]==0);

                                                            assert property (coverage0[175]==0);

                                                            assert property (coverage0[177]==0);

                                                            assert property (coverage0[181]==0);

                                                            assert property (coverage0[185]==0);

                                                    assert property (coverage0[191]==0);

                                                            assert property (coverage0[192]==0);

                                                            assert property (coverage0[194]==0);

                                                            assert property (coverage0[198]==0);

                                                            assert property (coverage0[202]==0);

                                                            assert property (coverage0[206]==0);

                                                            assert property (coverage0[208]==0);

                                                            assert property (coverage0[210]==0);

                                                            assert property (coverage0[212]==0);

                                                    assert property (coverage0[214]==0);

                                                            assert property (coverage0[215]==0);

                                                            assert property (coverage0[217]==0);

                                                            assert property (coverage0[221]==0);

                                                            assert property (coverage0[225]==0);

                                                            assert property (coverage0[229]==0);

                                                            assert property (coverage0[231]==0);

                                                            assert property (coverage0[233]==0);

                                                            assert property (coverage0[235]==0);

                                                    assert property (coverage0[237]==0);

                                                            assert property (coverage0[238]==0);

                                                            assert property (coverage0[240]==0);

                                                            assert property (coverage0[244]==0);

                                                            assert property (coverage0[248]==0);

                                                            assert property (coverage0[252]==0);

                                                            assert property (coverage0[254]==0);

                                                            assert property (coverage0[256]==0);

                                                            assert property (coverage0[258]==0);

                                                    assert property (coverage0[260]==0);

                                                            assert property (coverage0[261]==0);

                                                            assert property (coverage0[263]==0);

                                                            assert property (coverage0[267]==0);

                                                            assert property (coverage0[271]==0);

                                                            assert property (coverage0[275]==0);

                                                            assert property (coverage0[277]==0);

                                                            assert property (coverage0[279]==0);

                                                            assert property (coverage0[281]==0);

                                                    assert property (coverage0[283]==0);

                                                            assert property (coverage0[284]==0);

                                                            assert property (coverage0[286]==0);

                                                            assert property (coverage0[290]==0);

                                                            assert property (coverage0[294]==0);

                                                            assert property (coverage0[298]==0);

                                                            assert property (coverage0[300]==0);

                                                            assert property (coverage0[302]==0);

                                                            assert property (coverage0[304]==0);

                                                    assert property (coverage0[306]==0);

                                                            assert property (coverage0[307]==0);

                                                            assert property (coverage0[309]==0);

                                                            assert property (coverage0[313]==0);

                                                            assert property (coverage0[317]==0);

                                                            assert property (coverage0[321]==0);

                                                            assert property (coverage0[323]==0);

                                                            assert property (coverage0[325]==0);

                                                            assert property (coverage0[327]==0);

                                                    assert property (coverage0[329]==0);

                                                            assert property (coverage0[330]==0);

                                                            assert property (coverage0[332]==0);

                                                            assert property (coverage0[336]==0);

                                                            assert property (coverage0[340]==0);

                                                            assert property (coverage0[344]==0);

                                                            assert property (coverage0[346]==0);

                                                            assert property (coverage0[348]==0);

                                                            assert property (coverage0[350]==0);

                                                    assert property (coverage0[352]==0);

                                                            assert property (coverage0[353]==0);

                                                            assert property (coverage0[355]==0);

                                                            assert property (coverage0[359]==0);

                                                            assert property (coverage0[363]==0);

                                                            assert property (coverage0[367]==0);

                                                            assert property (coverage0[369]==0);

                                                            assert property (coverage0[371]==0);

                                                            assert property (coverage0[373]==0);

                                                    assert property (coverage0[375]==0);

                                                            assert property (coverage0[376]==0);

                                                            assert property (coverage0[378]==0);

                                                            assert property (coverage0[382]==0);

                                                            assert property (coverage0[386]==0);

                                                            assert property (coverage0[390]==0);

                                                            assert property (coverage0[392]==0);

                                                            assert property (coverage0[394]==0);

                                                            assert property (coverage0[396]==0);

                                                    assert property (coverage0[398]==0);

                                                            assert property (coverage0[399]==0);

                                                            assert property (coverage0[401]==0);

                                                            assert property (coverage0[405]==0);

                                                            assert property (coverage0[409]==0);

                                                            assert property (coverage0[413]==0);

                                                            assert property (coverage0[415]==0);

                                                            assert property (coverage0[417]==0);

                                                            assert property (coverage0[419]==0);

                                                    assert property (coverage0[421]==0);

                                                            assert property (coverage0[422]==0);

                                                            assert property (coverage0[424]==0);

                                                            assert property (coverage0[426]==0);

                                                            assert property (coverage0[428]==0);

                                                                    assert property (coverage0[430]==0);

                                                                    assert property (coverage0[431]==0);

                                                            assert property (coverage0[434]==0);

                                                            assert property (coverage0[436]==0);

                                                            assert property (coverage0[438]==0);

                                                            assert property (coverage0[440]==0);

                                            assert property (coverage0[145]==0);

                                                    assert property (coverage0[442]==0);

                                                            assert property (coverage0[444]==0);

                                                            assert property (coverage0[446]==0);

                                                            assert property (coverage0[448]==0);

                                                            assert property (coverage0[450]==0);

                                                    assert property (coverage0[443]==0);

endmodule
